
module processor (
	clk_clk,
	my_register_slave_interface_0_conduit_end_readdata,
	uart_0_rxd,
	uart_0_txd);	

	input		clk_clk;
	output	[31:0]	my_register_slave_interface_0_conduit_end_readdata;
	input		uart_0_rxd;
	output		uart_0_txd;
endmodule
